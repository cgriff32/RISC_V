// imem.v

// Generated using ACDS version 13.0 156 at 2019.07.16.14:23:04

`timescale 1 ps / 1 ps
module chip_mem (
		input  wire        clk_clk,             //     clk.clk
		input  wire        reset_reset_n,       //   reset.reset_n
		input  wire [9:0]  imem_in_address,     // imem_in.address
		input  wire        imem_in_debugaccess, //        .debugaccess
		input  wire        imem_in_clken,       //        .clken
		input  wire        imem_in_chipselect,  //        .chipselect
		input  wire        imem_in_write,       //        .write
		output wire [31:0] imem_in_readdata,    //        .readdata
		input  wire [31:0] imem_in_writedata,   //        .writedata
		input  wire [3:0]  imem_in_byteenable,  //        .byteenable
		input  wire [11:0] dmem_in_address,     // dmem_in.address
		input  wire        dmem_in_clken,       //        .clken
		input  wire        dmem_in_chipselect,  //        .chipselect
		input  wire        dmem_in_write,       //        .write
		output wire [7:0]  dmem_in_readdata,    //        .readdata
		input  wire [7:0]  dmem_in_writedata    //        .writedata
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> [dmem:reset, imem:reset]

	imem_imem imem (
		.clk         (clk_clk),                        //   clk1.clk
		.address     (imem_in_address),                //     s1.address
		.debugaccess (imem_in_debugaccess),            //       .debugaccess
		.clken       (imem_in_clken),                  //       .clken
		.chipselect  (imem_in_chipselect),             //       .chipselect
		.write       (imem_in_write),                  //       .write
		.readdata    (imem_in_readdata),               //       .readdata
		.writedata   (imem_in_writedata),              //       .writedata
		.byteenable  (imem_in_byteenable),             //       .byteenable
		.reset       (rst_controller_reset_out_reset)  // reset1.reset
	);

	imem_dmem dmem (
		.clk        (clk_clk),                        //   clk1.clk
		.address    (dmem_in_address),                //     s1.address
		.clken      (dmem_in_clken),                  //       .clken
		.chipselect (dmem_in_chipselect),             //       .chipselect
		.write      (dmem_in_write),                  //       .write
		.readdata   (dmem_in_readdata),               //       .readdata
		.writedata  (dmem_in_writedata),              //       .writedata
		.reset      (rst_controller_reset_out_reset)  // reset1.reset
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule

//
`include "constants.vh"